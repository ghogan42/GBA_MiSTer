module gba_colors
(
	input		enable,
	input		[7:0]	r, g, b,
	output	[7:0] r_out, g_out, b_out
);

wire	[9:0]	r_lin, g_lin, b_lin;
wire	[9:0]	r_gba, g_gba, b_gba;
wire	[7:0]	r_gba2, g_gba2, b_gba2;


// Convert from srgb to linear. I'm using srgb and not gamma 2.2 because precision
// is better on srgb for dark colors.

// Note that the output is 10 bits per channel
	srgb_to_linear(r,r_lin);
	srgb_to_linear(g,g_lin);
	srgb_to_linear(b,b_lin);

	
	
	
// Bit-shifting approximate GBA Colors
// This actually looks fine but you still have to do gamma to be close to correct
//always @(*) begin
//	gba_r = lin_r[9:1] + lin_r[9:2] + lin_r[9:3] + lin_g[9:3];
//	gba_g = lin_g[9:1] + lin_g[9:3] + lin_r[9:3] + lin_b[9:2];
//	gba_b = lin_b[9:1] + lin_b[9:2] + lin_r[9:3] + lin_r[9:4] + lin_g[9:4];
//end




//Calculate "GBA COlors" using the color mixer formula from the pixel shader
//out_r = 0.860*r + 0.190*g - 0.05*b
//out_g = 0.110*r + 0.660*g + 0.230*b
//out_b = 0.1325*r + 0.0575*g + 0.810*b

wire [19:0]	r_signed, g_signed, b_signed;
always @(*) begin
	r_signed = r_lin*(10'd220) + g_lin*(10'd49)  - b_lin*(10'd13);
	g_signed = r_lin*(10'd28)  + g_lin*(10'd169) + b_lin*(10'd59);
	b_signed = r_lin*(10'd34)  + g_lin*(10'd15)  + b_lin*(10'd207);
end


//Hopefully this will saturate values to 0 and 1023
assign r_gba = r_signed[19] ? 10'd0 : (r_signed[18] ? 10'd1023 : r_signed[17:8]);
assign g_gba = g_signed[19] ? 10'd0 : (g_signed[18] ? 10'd1023 : g_signed[17:8]);
assign b_gba = b_signed[19] ? 10'd0 : (b_signed[18] ? 10'd1023 : b_signed[17:8]);


// Now convert back to srgb space.  Input is 10 bits per channel and output is 8 bits per channel
linear_to_srgb(r_gba, r_gba2);
linear_to_srgb(g_gba, g_gba2);
linear_to_srgb(b_gba, b_gba2);

//Only change colors when module is enabled
assign r_out = enable ? r_gba2 : r;
assign g_out = enable ? g_gba2 : g;
assign b_out = enable ? b_gba2 : b;

endmodule


module srgb_to_linear
(
	input		[7:0]	col,
	output	[9	:0] out_col
);


always @(*) begin
	case (col)
		8'd0  :  out_col <= 10'd0;
		8'd1  :  out_col <= 10'd0;
		8'd2  :  out_col <= 10'd1;
		8'd3  :  out_col <= 10'd1;
		8'd4  :  out_col <= 10'd1;
		8'd5  :  out_col <= 10'd2;
		8'd6  :  out_col <= 10'd2;
		8'd7  :  out_col <= 10'd2;
		8'd8  :  out_col <= 10'd2;
		8'd9  :  out_col <= 10'd3;
		8'd10  :  out_col <= 10'd3;
		8'd11  :  out_col <= 10'd3;
		8'd12  :  out_col <= 10'd4;
		8'd13  :  out_col <= 10'd4;
		8'd14  :  out_col <= 10'd4;
		8'd15  :  out_col <= 10'd5;
		8'd16  :  out_col <= 10'd5;
		8'd17  :  out_col <= 10'd6;
		8'd18  :  out_col <= 10'd6;
		8'd19  :  out_col <= 10'd7;
		8'd20  :  out_col <= 10'd7;
		8'd21  :  out_col <= 10'd8;
		8'd22  :  out_col <= 10'd8;
		8'd23  :  out_col <= 10'd9;
		8'd24  :  out_col <= 10'd9;
		8'd25  :  out_col <= 10'd10;
		8'd26  :  out_col <= 10'd11;
		8'd27  :  out_col <= 10'd11;
		8'd28  :  out_col <= 10'd12;
		8'd29  :  out_col <= 10'd13;
		8'd30  :  out_col <= 10'd13;
		8'd31  :  out_col <= 10'd14;
		8'd32  :  out_col <= 10'd15;
		8'd33  :  out_col <= 10'd16;
		8'd34  :  out_col <= 10'd16;
		8'd35  :  out_col <= 10'd17;
		8'd36  :  out_col <= 10'd18;
		8'd37  :  out_col <= 10'd19;
		8'd38  :  out_col <= 10'd20;
		8'd39  :  out_col <= 10'd21;
		8'd40  :  out_col <= 10'd22;
		8'd41  :  out_col <= 10'd23;
		8'd42  :  out_col <= 10'd24;
		8'd43  :  out_col <= 10'd25;
		8'd44  :  out_col <= 10'd26;
		8'd45  :  out_col <= 10'd27;
		8'd46  :  out_col <= 10'd28;
		8'd47  :  out_col <= 10'd29;
		8'd48  :  out_col <= 10'd30;
		8'd49  :  out_col <= 10'd31;
		8'd50  :  out_col <= 10'd33;
		8'd51  :  out_col <= 10'd34;
		8'd52  :  out_col <= 10'd35;
		8'd53  :  out_col <= 10'd36;
		8'd54  :  out_col <= 10'd38;
		8'd55  :  out_col <= 10'd39;
		8'd56  :  out_col <= 10'd40;
		8'd57  :  out_col <= 10'd42;
		8'd58  :  out_col <= 10'd43;
		8'd59  :  out_col <= 10'd45;
		8'd60  :  out_col <= 10'd46;
		8'd61  :  out_col <= 10'd48;
		8'd62  :  out_col <= 10'd49;
		8'd63  :  out_col <= 10'd51;
		8'd64  :  out_col <= 10'd52;
		8'd65  :  out_col <= 10'd54;
		8'd66  :  out_col <= 10'd56;
		8'd67  :  out_col <= 10'd57;
		8'd68  :  out_col <= 10'd59;
		8'd69  :  out_col <= 10'd61;
		8'd70  :  out_col <= 10'd63;
		8'd71  :  out_col <= 10'd64;
		8'd72  :  out_col <= 10'd66;
		8'd73  :  out_col <= 10'd68;
		8'd74  :  out_col <= 10'd70;
		8'd75  :  out_col <= 10'd72;
		8'd76  :  out_col <= 10'd74;
		8'd77  :  out_col <= 10'd76;
		8'd78  :  out_col <= 10'd78;
		8'd79  :  out_col <= 10'd80;
		8'd80  :  out_col <= 10'd82;
		8'd81  :  out_col <= 10'd84;
		8'd82  :  out_col <= 10'd86;
		8'd83  :  out_col <= 10'd88;
		8'd84  :  out_col <= 10'd91;
		8'd85  :  out_col <= 10'd93;
		8'd86  :  out_col <= 10'd95;
		8'd87  :  out_col <= 10'd97;
		8'd88  :  out_col <= 10'd100;
		8'd89  :  out_col <= 10'd102;
		8'd90  :  out_col <= 10'd105;
		8'd91  :  out_col <= 10'd107;
		8'd92  :  out_col <= 10'd109;
		8'd93  :  out_col <= 10'd112;
		8'd94  :  out_col <= 10'd115;
		8'd95  :  out_col <= 10'd117;
		8'd96  :  out_col <= 10'd120;
		8'd97  :  out_col <= 10'd122;
		8'd98  :  out_col <= 10'd125;
		8'd99  :  out_col <= 10'd128;
		8'd100  :  out_col <= 10'd130;
		8'd101  :  out_col <= 10'd133;
		8'd102  :  out_col <= 10'd136;
		8'd103  :  out_col <= 10'd139;
		8'd104  :  out_col <= 10'd142;
		8'd105  :  out_col <= 10'd145;
		8'd106  :  out_col <= 10'd147;
		8'd107  :  out_col <= 10'd150;
		8'd108  :  out_col <= 10'd153;
		8'd109  :  out_col <= 10'd156;
		8'd110  :  out_col <= 10'd160;
		8'd111  :  out_col <= 10'd163;
		8'd112  :  out_col <= 10'd166;
		8'd113  :  out_col <= 10'd169;
		8'd114  :  out_col <= 10'd172;
		8'd115  :  out_col <= 10'd175;
		8'd116  :  out_col <= 10'd179;
		8'd117  :  out_col <= 10'd182;
		8'd118  :  out_col <= 10'd185;
		8'd119  :  out_col <= 10'd189;
		8'd120  :  out_col <= 10'd192;
		8'd121  :  out_col <= 10'd196;
		8'd122  :  out_col <= 10'd199;
		8'd123  :  out_col <= 10'd203;
		8'd124  :  out_col <= 10'd206;
		8'd125  :  out_col <= 10'd210;
		8'd126  :  out_col <= 10'd213;
		8'd127  :  out_col <= 10'd217;
		8'd128  :  out_col <= 10'd221;
		8'd129  :  out_col <= 10'd225;
		8'd130  :  out_col <= 10'd228;
		8'd131  :  out_col <= 10'd232;
		8'd132  :  out_col <= 10'd236;
		8'd133  :  out_col <= 10'd240;
		8'd134  :  out_col <= 10'd244;
		8'd135  :  out_col <= 10'd248;
		8'd136  :  out_col <= 10'd252;
		8'd137  :  out_col <= 10'd256;
		8'd138  :  out_col <= 10'd260;
		8'd139  :  out_col <= 10'd264;
		8'd140  :  out_col <= 10'd268;
		8'd141  :  out_col <= 10'd272;
		8'd142  :  out_col <= 10'd277;
		8'd143  :  out_col <= 10'd281;
		8'd144  :  out_col <= 10'd285;
		8'd145  :  out_col <= 10'd290;
		8'd146  :  out_col <= 10'd294;
		8'd147  :  out_col <= 10'd298;
		8'd148  :  out_col <= 10'd303;
		8'd149  :  out_col <= 10'd307;
		8'd150  :  out_col <= 10'd312;
		8'd151  :  out_col <= 10'd317;
		8'd152  :  out_col <= 10'd321;
		8'd153  :  out_col <= 10'd326;
		8'd154  :  out_col <= 10'd331;
		8'd155  :  out_col <= 10'd335;
		8'd156  :  out_col <= 10'd340;
		8'd157  :  out_col <= 10'd345;
		8'd158  :  out_col <= 10'd350;
		8'd159  :  out_col <= 10'd355;
		8'd160  :  out_col <= 10'd360;
		8'd161  :  out_col <= 10'd365;
		8'd162  :  out_col <= 10'd370;
		8'd163  :  out_col <= 10'd375;
		8'd164  :  out_col <= 10'd380;
		8'd165  :  out_col <= 10'd385;
		8'd166  :  out_col <= 10'd390;
		8'd167  :  out_col <= 10'd395;
		8'd168  :  out_col <= 10'd401;
		8'd169  :  out_col <= 10'd406;
		8'd170  :  out_col <= 10'd411;
		8'd171  :  out_col <= 10'd417;
		8'd172  :  out_col <= 10'd422;
		8'd173  :  out_col <= 10'd427;
		8'd174  :  out_col <= 10'd433;
		8'd175  :  out_col <= 10'd439;
		8'd176  :  out_col <= 10'd444;
		8'd177  :  out_col <= 10'd450;
		8'd178  :  out_col <= 10'd455;
		8'd179  :  out_col <= 10'd461;
		8'd180  :  out_col <= 10'd467;
		8'd181  :  out_col <= 10'd473;
		8'd182  :  out_col <= 10'd479;
		8'd183  :  out_col <= 10'd484;
		8'd184  :  out_col <= 10'd490;
		8'd185  :  out_col <= 10'd496;
		8'd186  :  out_col <= 10'd502;
		8'd187  :  out_col <= 10'd508;
		8'd188  :  out_col <= 10'd514;
		8'd189  :  out_col <= 10'd521;
		8'd190  :  out_col <= 10'd527;
		8'd191  :  out_col <= 10'd533;
		8'd192  :  out_col <= 10'd539;
		8'd193  :  out_col <= 10'd546;
		8'd194  :  out_col <= 10'd552;
		8'd195  :  out_col <= 10'd558;
		8'd196  :  out_col <= 10'd565;
		8'd197  :  out_col <= 10'd571;
		8'd198  :  out_col <= 10'd578;
		8'd199  :  out_col <= 10'd584;
		8'd200  :  out_col <= 10'd591;
		8'd201  :  out_col <= 10'd598;
		8'd202  :  out_col <= 10'd604;
		8'd203  :  out_col <= 10'd611;
		8'd204  :  out_col <= 10'd618;
		8'd205  :  out_col <= 10'd625;
		8'd206  :  out_col <= 10'd631;
		8'd207  :  out_col <= 10'd638;
		8'd208  :  out_col <= 10'd645;
		8'd209  :  out_col <= 10'd652;
		8'd210  :  out_col <= 10'd659;
		8'd211  :  out_col <= 10'd666;
		8'd212  :  out_col <= 10'd674;
		8'd213  :  out_col <= 10'd681;
		8'd214  :  out_col <= 10'd688;
		8'd215  :  out_col <= 10'd695;
		8'd216  :  out_col <= 10'd702;
		8'd217  :  out_col <= 10'd710;
		8'd218  :  out_col <= 10'd717;
		8'd219  :  out_col <= 10'd725;
		8'd220  :  out_col <= 10'd732;
		8'd221  :  out_col <= 10'd740;
		8'd222  :  out_col <= 10'd747;
		8'd223  :  out_col <= 10'd755;
		8'd224  :  out_col <= 10'd763;
		8'd225  :  out_col <= 10'd770;
		8'd226  :  out_col <= 10'd778;
		8'd227  :  out_col <= 10'd786;
		8'd228  :  out_col <= 10'd794;
		8'd229  :  out_col <= 10'd802;
		8'd230  :  out_col <= 10'd809;
		8'd231  :  out_col <= 10'd817;
		8'd232  :  out_col <= 10'd826;
		8'd233  :  out_col <= 10'd834;
		8'd234  :  out_col <= 10'd842;
		8'd235  :  out_col <= 10'd850;
		8'd236  :  out_col <= 10'd858;
		8'd237  :  out_col <= 10'd866;
		8'd238  :  out_col <= 10'd875;
		8'd239  :  out_col <= 10'd883;
		8'd240  :  out_col <= 10'd891;
		8'd241  :  out_col <= 10'd900;
		8'd242  :  out_col <= 10'd908;
		8'd243  :  out_col <= 10'd917;
		8'd244  :  out_col <= 10'd925;
		8'd245  :  out_col <= 10'd934;
		8'd246  :  out_col <= 10'd943;
		8'd247  :  out_col <= 10'd952;
		8'd248  :  out_col <= 10'd960;
		8'd249  :  out_col <= 10'd969;
		8'd250  :  out_col <= 10'd978;
		8'd251  :  out_col <= 10'd987;
		8'd252  :  out_col <= 10'd996;
		8'd253  :  out_col <= 10'd1005;
		8'd254  :  out_col <= 10'd1014;
		8'd255  :  out_col <= 10'd1023;
		default :  out_col <= 10'd0;
	endcase
end
endmodule


//linear to srgb uses a 10 bit table.  That's still not enough for full precision...
module linear_to_srgb
(
	input		[9:0]	col,
	output	[7:0] out_col
);


always @(*) begin
	case (col)
		10'd0  :  out_col <= 8'd0;
		10'd1  :  out_col <= 8'd3;
		10'd2  :  out_col <= 8'd6;
		10'd3  :  out_col <= 8'd10;
		10'd4  :  out_col <= 8'd13;
		10'd5  :  out_col <= 8'd15;
		10'd6  :  out_col <= 8'd18;
		10'd7  :  out_col <= 8'd20;
		10'd8  :  out_col <= 8'd22;
		10'd9  :  out_col <= 8'd23;
		10'd10  :  out_col <= 8'd25;
		10'd11  :  out_col <= 8'd27;
		10'd12  :  out_col <= 8'd28;
		10'd13  :  out_col <= 8'd30;
		10'd14  :  out_col <= 8'd31;
		10'd15  :  out_col <= 8'd32;
		10'd16  :  out_col <= 8'd34;
		10'd17  :  out_col <= 8'd35;
		10'd18  :  out_col <= 8'd36;
		10'd19  :  out_col <= 8'd37;
		10'd20  :  out_col <= 8'd38;
		10'd21  :  out_col <= 8'd39;
		10'd22  :  out_col <= 8'd40;
		10'd23  :  out_col <= 8'd41;
		10'd24  :  out_col <= 8'd42;
		10'd25  :  out_col <= 8'd43;
		10'd26  :  out_col <= 8'd44;
		10'd27  :  out_col <= 8'd45;
		10'd28  :  out_col <= 8'd46;
		10'd29  :  out_col <= 8'd47;
		10'd30  :  out_col <= 8'd48;
		10'd31  :  out_col <= 8'd49;
		10'd32  :  out_col <= 8'd49;
		10'd33  :  out_col <= 8'd50;
		10'd34  :  out_col <= 8'd51;
		10'd35  :  out_col <= 8'd52;
		10'd36  :  out_col <= 8'd53;
		10'd37  :  out_col <= 8'd53;
		10'd38  :  out_col <= 8'd54;
		10'd39  :  out_col <= 8'd55;
		10'd40  :  out_col <= 8'd56;
		10'd41  :  out_col <= 8'd56;
		10'd42  :  out_col <= 8'd57;
		10'd43  :  out_col <= 8'd58;
		10'd44  :  out_col <= 8'd58;
		10'd45  :  out_col <= 8'd59;
		10'd46  :  out_col <= 8'd60;
		10'd47  :  out_col <= 8'd61;
		10'd48  :  out_col <= 8'd61;
		10'd49  :  out_col <= 8'd62;
		10'd50  :  out_col <= 8'd62;
		10'd51  :  out_col <= 8'd63;
		10'd52  :  out_col <= 8'd64;
		10'd53  :  out_col <= 8'd64;
		10'd54  :  out_col <= 8'd65;
		10'd55  :  out_col <= 8'd66;
		10'd56  :  out_col <= 8'd66;
		10'd57  :  out_col <= 8'd67;
		10'd58  :  out_col <= 8'd67;
		10'd59  :  out_col <= 8'd68;
		10'd60  :  out_col <= 8'd68;
		10'd61  :  out_col <= 8'd69;
		10'd62  :  out_col <= 8'd70;
		10'd63  :  out_col <= 8'd70;
		10'd64  :  out_col <= 8'd71;
		10'd65  :  out_col <= 8'd71;
		10'd66  :  out_col <= 8'd72;
		10'd67  :  out_col <= 8'd72;
		10'd68  :  out_col <= 8'd73;
		10'd69  :  out_col <= 8'd73;
		10'd70  :  out_col <= 8'd74;
		10'd71  :  out_col <= 8'd74;
		10'd72  :  out_col <= 8'd75;
		10'd73  :  out_col <= 8'd76;
		10'd74  :  out_col <= 8'd76;
		10'd75  :  out_col <= 8'd77;
		10'd76  :  out_col <= 8'd77;
		10'd77  :  out_col <= 8'd78;
		10'd78  :  out_col <= 8'd78;
		10'd79  :  out_col <= 8'd79;
		10'd80  :  out_col <= 8'd79;
		10'd81  :  out_col <= 8'd79;
		10'd82  :  out_col <= 8'd80;
		10'd83  :  out_col <= 8'd80;
		10'd84  :  out_col <= 8'd81;
		10'd85  :  out_col <= 8'd81;
		10'd86  :  out_col <= 8'd82;
		10'd87  :  out_col <= 8'd82;
		10'd88  :  out_col <= 8'd83;
		10'd89  :  out_col <= 8'd83;
		10'd90  :  out_col <= 8'd84;
		10'd91  :  out_col <= 8'd84;
		10'd92  :  out_col <= 8'd85;
		10'd93  :  out_col <= 8'd85;
		10'd94  :  out_col <= 8'd85;
		10'd95  :  out_col <= 8'd86;
		10'd96  :  out_col <= 8'd86;
		10'd97  :  out_col <= 8'd87;
		10'd98  :  out_col <= 8'd87;
		10'd99  :  out_col <= 8'd88;
		10'd100  :  out_col <= 8'd88;
		10'd101  :  out_col <= 8'd88;
		10'd102  :  out_col <= 8'd89;
		10'd103  :  out_col <= 8'd89;
		10'd104  :  out_col <= 8'd90;
		10'd105  :  out_col <= 8'd90;
		10'd106  :  out_col <= 8'd91;
		10'd107  :  out_col <= 8'd91;
		10'd108  :  out_col <= 8'd91;
		10'd109  :  out_col <= 8'd92;
		10'd110  :  out_col <= 8'd92;
		10'd111  :  out_col <= 8'd93;
		10'd112  :  out_col <= 8'd93;
		10'd113  :  out_col <= 8'd93;
		10'd114  :  out_col <= 8'd94;
		10'd115  :  out_col <= 8'd94;
		10'd116  :  out_col <= 8'd95;
		10'd117  :  out_col <= 8'd95;
		10'd118  :  out_col <= 8'd95;
		10'd119  :  out_col <= 8'd96;
		10'd120  :  out_col <= 8'd96;
		10'd121  :  out_col <= 8'd97;
		10'd122  :  out_col <= 8'd97;
		10'd123  :  out_col <= 8'd97;
		10'd124  :  out_col <= 8'd98;
		10'd125  :  out_col <= 8'd98;
		10'd126  :  out_col <= 8'd98;
		10'd127  :  out_col <= 8'd99;
		10'd128  :  out_col <= 8'd99;
		10'd129  :  out_col <= 8'd99;
		10'd130  :  out_col <= 8'd100;
		10'd131  :  out_col <= 8'd100;
		10'd132  :  out_col <= 8'd101;
		10'd133  :  out_col <= 8'd101;
		10'd134  :  out_col <= 8'd101;
		10'd135  :  out_col <= 8'd102;
		10'd136  :  out_col <= 8'd102;
		10'd137  :  out_col <= 8'd102;
		10'd138  :  out_col <= 8'd103;
		10'd139  :  out_col <= 8'd103;
		10'd140  :  out_col <= 8'd103;
		10'd141  :  out_col <= 8'd104;
		10'd142  :  out_col <= 8'd104;
		10'd143  :  out_col <= 8'd104;
		10'd144  :  out_col <= 8'd105;
		10'd145  :  out_col <= 8'd105;
		10'd146  :  out_col <= 8'd106;
		10'd147  :  out_col <= 8'd106;
		10'd148  :  out_col <= 8'd106;
		10'd149  :  out_col <= 8'd107;
		10'd150  :  out_col <= 8'd107;
		10'd151  :  out_col <= 8'd107;
		10'd152  :  out_col <= 8'd108;
		10'd153  :  out_col <= 8'd108;
		10'd154  :  out_col <= 8'd108;
		10'd155  :  out_col <= 8'd109;
		10'd156  :  out_col <= 8'd109;
		10'd157  :  out_col <= 8'd109;
		10'd158  :  out_col <= 8'd110;
		10'd159  :  out_col <= 8'd110;
		10'd160  :  out_col <= 8'd110;
		10'd161  :  out_col <= 8'd110;
		10'd162  :  out_col <= 8'd111;
		10'd163  :  out_col <= 8'd111;
		10'd164  :  out_col <= 8'd111;
		10'd165  :  out_col <= 8'd112;
		10'd166  :  out_col <= 8'd112;
		10'd167  :  out_col <= 8'd112;
		10'd168  :  out_col <= 8'd113;
		10'd169  :  out_col <= 8'd113;
		10'd170  :  out_col <= 8'd113;
		10'd171  :  out_col <= 8'd114;
		10'd172  :  out_col <= 8'd114;
		10'd173  :  out_col <= 8'd114;
		10'd174  :  out_col <= 8'd115;
		10'd175  :  out_col <= 8'd115;
		10'd176  :  out_col <= 8'd115;
		10'd177  :  out_col <= 8'd115;
		10'd178  :  out_col <= 8'd116;
		10'd179  :  out_col <= 8'd116;
		10'd180  :  out_col <= 8'd116;
		10'd181  :  out_col <= 8'd117;
		10'd182  :  out_col <= 8'd117;
		10'd183  :  out_col <= 8'd117;
		10'd184  :  out_col <= 8'd118;
		10'd185  :  out_col <= 8'd118;
		10'd186  :  out_col <= 8'd118;
		10'd187  :  out_col <= 8'd118;
		10'd188  :  out_col <= 8'd119;
		10'd189  :  out_col <= 8'd119;
		10'd190  :  out_col <= 8'd119;
		10'd191  :  out_col <= 8'd120;
		10'd192  :  out_col <= 8'd120;
		10'd193  :  out_col <= 8'd120;
		10'd194  :  out_col <= 8'd121;
		10'd195  :  out_col <= 8'd121;
		10'd196  :  out_col <= 8'd121;
		10'd197  :  out_col <= 8'd121;
		10'd198  :  out_col <= 8'd122;
		10'd199  :  out_col <= 8'd122;
		10'd200  :  out_col <= 8'd122;
		10'd201  :  out_col <= 8'd123;
		10'd202  :  out_col <= 8'd123;
		10'd203  :  out_col <= 8'd123;
		10'd204  :  out_col <= 8'd123;
		10'd205  :  out_col <= 8'd124;
		10'd206  :  out_col <= 8'd124;
		10'd207  :  out_col <= 8'd124;
		10'd208  :  out_col <= 8'd125;
		10'd209  :  out_col <= 8'd125;
		10'd210  :  out_col <= 8'd125;
		10'd211  :  out_col <= 8'd125;
		10'd212  :  out_col <= 8'd126;
		10'd213  :  out_col <= 8'd126;
		10'd214  :  out_col <= 8'd126;
		10'd215  :  out_col <= 8'd126;
		10'd216  :  out_col <= 8'd127;
		10'd217  :  out_col <= 8'd127;
		10'd218  :  out_col <= 8'd127;
		10'd219  :  out_col <= 8'd128;
		10'd220  :  out_col <= 8'd128;
		10'd221  :  out_col <= 8'd128;
		10'd222  :  out_col <= 8'd128;
		10'd223  :  out_col <= 8'd129;
		10'd224  :  out_col <= 8'd129;
		10'd225  :  out_col <= 8'd129;
		10'd226  :  out_col <= 8'd129;
		10'd227  :  out_col <= 8'd130;
		10'd228  :  out_col <= 8'd130;
		10'd229  :  out_col <= 8'd130;
		10'd230  :  out_col <= 8'd130;
		10'd231  :  out_col <= 8'd131;
		10'd232  :  out_col <= 8'd131;
		10'd233  :  out_col <= 8'd131;
		10'd234  :  out_col <= 8'd131;
		10'd235  :  out_col <= 8'd132;
		10'd236  :  out_col <= 8'd132;
		10'd237  :  out_col <= 8'd132;
		10'd238  :  out_col <= 8'd133;
		10'd239  :  out_col <= 8'd133;
		10'd240  :  out_col <= 8'd133;
		10'd241  :  out_col <= 8'd133;
		10'd242  :  out_col <= 8'd134;
		10'd243  :  out_col <= 8'd134;
		10'd244  :  out_col <= 8'd134;
		10'd245  :  out_col <= 8'd134;
		10'd246  :  out_col <= 8'd135;
		10'd247  :  out_col <= 8'd135;
		10'd248  :  out_col <= 8'd135;
		10'd249  :  out_col <= 8'd135;
		10'd250  :  out_col <= 8'd136;
		10'd251  :  out_col <= 8'd136;
		10'd252  :  out_col <= 8'd136;
		10'd253  :  out_col <= 8'd136;
		10'd254  :  out_col <= 8'd137;
		10'd255  :  out_col <= 8'd137;
		10'd256  :  out_col <= 8'd137;
		10'd257  :  out_col <= 8'd137;
		10'd258  :  out_col <= 8'd138;
		10'd259  :  out_col <= 8'd138;
		10'd260  :  out_col <= 8'd138;
		10'd261  :  out_col <= 8'd138;
		10'd262  :  out_col <= 8'd138;
		10'd263  :  out_col <= 8'd139;
		10'd264  :  out_col <= 8'd139;
		10'd265  :  out_col <= 8'd139;
		10'd266  :  out_col <= 8'd139;
		10'd267  :  out_col <= 8'd140;
		10'd268  :  out_col <= 8'd140;
		10'd269  :  out_col <= 8'd140;
		10'd270  :  out_col <= 8'd140;
		10'd271  :  out_col <= 8'd141;
		10'd272  :  out_col <= 8'd141;
		10'd273  :  out_col <= 8'd141;
		10'd274  :  out_col <= 8'd141;
		10'd275  :  out_col <= 8'd142;
		10'd276  :  out_col <= 8'd142;
		10'd277  :  out_col <= 8'd142;
		10'd278  :  out_col <= 8'd142;
		10'd279  :  out_col <= 8'd143;
		10'd280  :  out_col <= 8'd143;
		10'd281  :  out_col <= 8'd143;
		10'd282  :  out_col <= 8'd143;
		10'd283  :  out_col <= 8'd143;
		10'd284  :  out_col <= 8'd144;
		10'd285  :  out_col <= 8'd144;
		10'd286  :  out_col <= 8'd144;
		10'd287  :  out_col <= 8'd144;
		10'd288  :  out_col <= 8'd145;
		10'd289  :  out_col <= 8'd145;
		10'd290  :  out_col <= 8'd145;
		10'd291  :  out_col <= 8'd145;
		10'd292  :  out_col <= 8'd146;
		10'd293  :  out_col <= 8'd146;
		10'd294  :  out_col <= 8'd146;
		10'd295  :  out_col <= 8'd146;
		10'd296  :  out_col <= 8'd146;
		10'd297  :  out_col <= 8'd147;
		10'd298  :  out_col <= 8'd147;
		10'd299  :  out_col <= 8'd147;
		10'd300  :  out_col <= 8'd147;
		10'd301  :  out_col <= 8'd148;
		10'd302  :  out_col <= 8'd148;
		10'd303  :  out_col <= 8'd148;
		10'd304  :  out_col <= 8'd148;
		10'd305  :  out_col <= 8'd148;
		10'd306  :  out_col <= 8'd149;
		10'd307  :  out_col <= 8'd149;
		10'd308  :  out_col <= 8'd149;
		10'd309  :  out_col <= 8'd149;
		10'd310  :  out_col <= 8'd150;
		10'd311  :  out_col <= 8'd150;
		10'd312  :  out_col <= 8'd150;
		10'd313  :  out_col <= 8'd150;
		10'd314  :  out_col <= 8'd150;
		10'd315  :  out_col <= 8'd151;
		10'd316  :  out_col <= 8'd151;
		10'd317  :  out_col <= 8'd151;
		10'd318  :  out_col <= 8'd151;
		10'd319  :  out_col <= 8'd152;
		10'd320  :  out_col <= 8'd152;
		10'd321  :  out_col <= 8'd152;
		10'd322  :  out_col <= 8'd152;
		10'd323  :  out_col <= 8'd152;
		10'd324  :  out_col <= 8'd153;
		10'd325  :  out_col <= 8'd153;
		10'd326  :  out_col <= 8'd153;
		10'd327  :  out_col <= 8'd153;
		10'd328  :  out_col <= 8'd153;
		10'd329  :  out_col <= 8'd154;
		10'd330  :  out_col <= 8'd154;
		10'd331  :  out_col <= 8'd154;
		10'd332  :  out_col <= 8'd154;
		10'd333  :  out_col <= 8'd155;
		10'd334  :  out_col <= 8'd155;
		10'd335  :  out_col <= 8'd155;
		10'd336  :  out_col <= 8'd155;
		10'd337  :  out_col <= 8'd155;
		10'd338  :  out_col <= 8'd156;
		10'd339  :  out_col <= 8'd156;
		10'd340  :  out_col <= 8'd156;
		10'd341  :  out_col <= 8'd156;
		10'd342  :  out_col <= 8'd156;
		10'd343  :  out_col <= 8'd157;
		10'd344  :  out_col <= 8'd157;
		10'd345  :  out_col <= 8'd157;
		10'd346  :  out_col <= 8'd157;
		10'd347  :  out_col <= 8'd157;
		10'd348  :  out_col <= 8'd158;
		10'd349  :  out_col <= 8'd158;
		10'd350  :  out_col <= 8'd158;
		10'd351  :  out_col <= 8'd158;
		10'd352  :  out_col <= 8'd158;
		10'd353  :  out_col <= 8'd159;
		10'd354  :  out_col <= 8'd159;
		10'd355  :  out_col <= 8'd159;
		10'd356  :  out_col <= 8'd159;
		10'd357  :  out_col <= 8'd159;
		10'd358  :  out_col <= 8'd160;
		10'd359  :  out_col <= 8'd160;
		10'd360  :  out_col <= 8'd160;
		10'd361  :  out_col <= 8'd160;
		10'd362  :  out_col <= 8'd160;
		10'd363  :  out_col <= 8'd161;
		10'd364  :  out_col <= 8'd161;
		10'd365  :  out_col <= 8'd161;
		10'd366  :  out_col <= 8'd161;
		10'd367  :  out_col <= 8'd161;
		10'd368  :  out_col <= 8'd162;
		10'd369  :  out_col <= 8'd162;
		10'd370  :  out_col <= 8'd162;
		10'd371  :  out_col <= 8'd162;
		10'd372  :  out_col <= 8'd162;
		10'd373  :  out_col <= 8'd163;
		10'd374  :  out_col <= 8'd163;
		10'd375  :  out_col <= 8'd163;
		10'd376  :  out_col <= 8'd163;
		10'd377  :  out_col <= 8'd163;
		10'd378  :  out_col <= 8'd164;
		10'd379  :  out_col <= 8'd164;
		10'd380  :  out_col <= 8'd164;
		10'd381  :  out_col <= 8'd164;
		10'd382  :  out_col <= 8'd164;
		10'd383  :  out_col <= 8'd165;
		10'd384  :  out_col <= 8'd165;
		10'd385  :  out_col <= 8'd165;
		10'd386  :  out_col <= 8'd165;
		10'd387  :  out_col <= 8'd165;
		10'd388  :  out_col <= 8'd166;
		10'd389  :  out_col <= 8'd166;
		10'd390  :  out_col <= 8'd166;
		10'd391  :  out_col <= 8'd166;
		10'd392  :  out_col <= 8'd166;
		10'd393  :  out_col <= 8'd167;
		10'd394  :  out_col <= 8'd167;
		10'd395  :  out_col <= 8'd167;
		10'd396  :  out_col <= 8'd167;
		10'd397  :  out_col <= 8'd167;
		10'd398  :  out_col <= 8'd168;
		10'd399  :  out_col <= 8'd168;
		10'd400  :  out_col <= 8'd168;
		10'd401  :  out_col <= 8'd168;
		10'd402  :  out_col <= 8'd168;
		10'd403  :  out_col <= 8'd168;
		10'd404  :  out_col <= 8'd169;
		10'd405  :  out_col <= 8'd169;
		10'd406  :  out_col <= 8'd169;
		10'd407  :  out_col <= 8'd169;
		10'd408  :  out_col <= 8'd169;
		10'd409  :  out_col <= 8'd170;
		10'd410  :  out_col <= 8'd170;
		10'd411  :  out_col <= 8'd170;
		10'd412  :  out_col <= 8'd170;
		10'd413  :  out_col <= 8'd170;
		10'd414  :  out_col <= 8'd171;
		10'd415  :  out_col <= 8'd171;
		10'd416  :  out_col <= 8'd171;
		10'd417  :  out_col <= 8'd171;
		10'd418  :  out_col <= 8'd171;
		10'd419  :  out_col <= 8'd171;
		10'd420  :  out_col <= 8'd172;
		10'd421  :  out_col <= 8'd172;
		10'd422  :  out_col <= 8'd172;
		10'd423  :  out_col <= 8'd172;
		10'd424  :  out_col <= 8'd172;
		10'd425  :  out_col <= 8'd173;
		10'd426  :  out_col <= 8'd173;
		10'd427  :  out_col <= 8'd173;
		10'd428  :  out_col <= 8'd173;
		10'd429  :  out_col <= 8'd173;
		10'd430  :  out_col <= 8'd173;
		10'd431  :  out_col <= 8'd174;
		10'd432  :  out_col <= 8'd174;
		10'd433  :  out_col <= 8'd174;
		10'd434  :  out_col <= 8'd174;
		10'd435  :  out_col <= 8'd174;
		10'd436  :  out_col <= 8'd175;
		10'd437  :  out_col <= 8'd175;
		10'd438  :  out_col <= 8'd175;
		10'd439  :  out_col <= 8'd175;
		10'd440  :  out_col <= 8'd175;
		10'd441  :  out_col <= 8'd175;
		10'd442  :  out_col <= 8'd176;
		10'd443  :  out_col <= 8'd176;
		10'd444  :  out_col <= 8'd176;
		10'd445  :  out_col <= 8'd176;
		10'd446  :  out_col <= 8'd176;
		10'd447  :  out_col <= 8'd177;
		10'd448  :  out_col <= 8'd177;
		10'd449  :  out_col <= 8'd177;
		10'd450  :  out_col <= 8'd177;
		10'd451  :  out_col <= 8'd177;
		10'd452  :  out_col <= 8'd177;
		10'd453  :  out_col <= 8'd178;
		10'd454  :  out_col <= 8'd178;
		10'd455  :  out_col <= 8'd178;
		10'd456  :  out_col <= 8'd178;
		10'd457  :  out_col <= 8'd178;
		10'd458  :  out_col <= 8'd178;
		10'd459  :  out_col <= 8'd179;
		10'd460  :  out_col <= 8'd179;
		10'd461  :  out_col <= 8'd179;
		10'd462  :  out_col <= 8'd179;
		10'd463  :  out_col <= 8'd179;
		10'd464  :  out_col <= 8'd179;
		10'd465  :  out_col <= 8'd180;
		10'd466  :  out_col <= 8'd180;
		10'd467  :  out_col <= 8'd180;
		10'd468  :  out_col <= 8'd180;
		10'd469  :  out_col <= 8'd180;
		10'd470  :  out_col <= 8'd181;
		10'd471  :  out_col <= 8'd181;
		10'd472  :  out_col <= 8'd181;
		10'd473  :  out_col <= 8'd181;
		10'd474  :  out_col <= 8'd181;
		10'd475  :  out_col <= 8'd181;
		10'd476  :  out_col <= 8'd182;
		10'd477  :  out_col <= 8'd182;
		10'd478  :  out_col <= 8'd182;
		10'd479  :  out_col <= 8'd182;
		10'd480  :  out_col <= 8'd182;
		10'd481  :  out_col <= 8'd182;
		10'd482  :  out_col <= 8'd183;
		10'd483  :  out_col <= 8'd183;
		10'd484  :  out_col <= 8'd183;
		10'd485  :  out_col <= 8'd183;
		10'd486  :  out_col <= 8'd183;
		10'd487  :  out_col <= 8'd183;
		10'd488  :  out_col <= 8'd184;
		10'd489  :  out_col <= 8'd184;
		10'd490  :  out_col <= 8'd184;
		10'd491  :  out_col <= 8'd184;
		10'd492  :  out_col <= 8'd184;
		10'd493  :  out_col <= 8'd184;
		10'd494  :  out_col <= 8'd185;
		10'd495  :  out_col <= 8'd185;
		10'd496  :  out_col <= 8'd185;
		10'd497  :  out_col <= 8'd185;
		10'd498  :  out_col <= 8'd185;
		10'd499  :  out_col <= 8'd185;
		10'd500  :  out_col <= 8'd186;
		10'd501  :  out_col <= 8'd186;
		10'd502  :  out_col <= 8'd186;
		10'd503  :  out_col <= 8'd186;
		10'd504  :  out_col <= 8'd186;
		10'd505  :  out_col <= 8'd186;
		10'd506  :  out_col <= 8'd187;
		10'd507  :  out_col <= 8'd187;
		10'd508  :  out_col <= 8'd187;
		10'd509  :  out_col <= 8'd187;
		10'd510  :  out_col <= 8'd187;
		10'd511  :  out_col <= 8'd187;
		10'd512  :  out_col <= 8'd188;
		10'd513  :  out_col <= 8'd188;
		10'd514  :  out_col <= 8'd188;
		10'd515  :  out_col <= 8'd188;
		10'd516  :  out_col <= 8'd188;
		10'd517  :  out_col <= 8'd188;
		10'd518  :  out_col <= 8'd189;
		10'd519  :  out_col <= 8'd189;
		10'd520  :  out_col <= 8'd189;
		10'd521  :  out_col <= 8'd189;
		10'd522  :  out_col <= 8'd189;
		10'd523  :  out_col <= 8'd189;
		10'd524  :  out_col <= 8'd190;
		10'd525  :  out_col <= 8'd190;
		10'd526  :  out_col <= 8'd190;
		10'd527  :  out_col <= 8'd190;
		10'd528  :  out_col <= 8'd190;
		10'd529  :  out_col <= 8'd190;
		10'd530  :  out_col <= 8'd191;
		10'd531  :  out_col <= 8'd191;
		10'd532  :  out_col <= 8'd191;
		10'd533  :  out_col <= 8'd191;
		10'd534  :  out_col <= 8'd191;
		10'd535  :  out_col <= 8'd191;
		10'd536  :  out_col <= 8'd191;
		10'd537  :  out_col <= 8'd192;
		10'd538  :  out_col <= 8'd192;
		10'd539  :  out_col <= 8'd192;
		10'd540  :  out_col <= 8'd192;
		10'd541  :  out_col <= 8'd192;
		10'd542  :  out_col <= 8'd192;
		10'd543  :  out_col <= 8'd193;
		10'd544  :  out_col <= 8'd193;
		10'd545  :  out_col <= 8'd193;
		10'd546  :  out_col <= 8'd193;
		10'd547  :  out_col <= 8'd193;
		10'd548  :  out_col <= 8'd193;
		10'd549  :  out_col <= 8'd194;
		10'd550  :  out_col <= 8'd194;
		10'd551  :  out_col <= 8'd194;
		10'd552  :  out_col <= 8'd194;
		10'd553  :  out_col <= 8'd194;
		10'd554  :  out_col <= 8'd194;
		10'd555  :  out_col <= 8'd194;
		10'd556  :  out_col <= 8'd195;
		10'd557  :  out_col <= 8'd195;
		10'd558  :  out_col <= 8'd195;
		10'd559  :  out_col <= 8'd195;
		10'd560  :  out_col <= 8'd195;
		10'd561  :  out_col <= 8'd195;
		10'd562  :  out_col <= 8'd196;
		10'd563  :  out_col <= 8'd196;
		10'd564  :  out_col <= 8'd196;
		10'd565  :  out_col <= 8'd196;
		10'd566  :  out_col <= 8'd196;
		10'd567  :  out_col <= 8'd196;
		10'd568  :  out_col <= 8'd197;
		10'd569  :  out_col <= 8'd197;
		10'd570  :  out_col <= 8'd197;
		10'd571  :  out_col <= 8'd197;
		10'd572  :  out_col <= 8'd197;
		10'd573  :  out_col <= 8'd197;
		10'd574  :  out_col <= 8'd197;
		10'd575  :  out_col <= 8'd198;
		10'd576  :  out_col <= 8'd198;
		10'd577  :  out_col <= 8'd198;
		10'd578  :  out_col <= 8'd198;
		10'd579  :  out_col <= 8'd198;
		10'd580  :  out_col <= 8'd198;
		10'd581  :  out_col <= 8'd199;
		10'd582  :  out_col <= 8'd199;
		10'd583  :  out_col <= 8'd199;
		10'd584  :  out_col <= 8'd199;
		10'd585  :  out_col <= 8'd199;
		10'd586  :  out_col <= 8'd199;
		10'd587  :  out_col <= 8'd199;
		10'd588  :  out_col <= 8'd200;
		10'd589  :  out_col <= 8'd200;
		10'd590  :  out_col <= 8'd200;
		10'd591  :  out_col <= 8'd200;
		10'd592  :  out_col <= 8'd200;
		10'd593  :  out_col <= 8'd200;
		10'd594  :  out_col <= 8'd200;
		10'd595  :  out_col <= 8'd201;
		10'd596  :  out_col <= 8'd201;
		10'd597  :  out_col <= 8'd201;
		10'd598  :  out_col <= 8'd201;
		10'd599  :  out_col <= 8'd201;
		10'd600  :  out_col <= 8'd201;
		10'd601  :  out_col <= 8'd202;
		10'd602  :  out_col <= 8'd202;
		10'd603  :  out_col <= 8'd202;
		10'd604  :  out_col <= 8'd202;
		10'd605  :  out_col <= 8'd202;
		10'd606  :  out_col <= 8'd202;
		10'd607  :  out_col <= 8'd202;
		10'd608  :  out_col <= 8'd203;
		10'd609  :  out_col <= 8'd203;
		10'd610  :  out_col <= 8'd203;
		10'd611  :  out_col <= 8'd203;
		10'd612  :  out_col <= 8'd203;
		10'd613  :  out_col <= 8'd203;
		10'd614  :  out_col <= 8'd203;
		10'd615  :  out_col <= 8'd204;
		10'd616  :  out_col <= 8'd204;
		10'd617  :  out_col <= 8'd204;
		10'd618  :  out_col <= 8'd204;
		10'd619  :  out_col <= 8'd204;
		10'd620  :  out_col <= 8'd204;
		10'd621  :  out_col <= 8'd204;
		10'd622  :  out_col <= 8'd205;
		10'd623  :  out_col <= 8'd205;
		10'd624  :  out_col <= 8'd205;
		10'd625  :  out_col <= 8'd205;
		10'd626  :  out_col <= 8'd205;
		10'd627  :  out_col <= 8'd205;
		10'd628  :  out_col <= 8'd206;
		10'd629  :  out_col <= 8'd206;
		10'd630  :  out_col <= 8'd206;
		10'd631  :  out_col <= 8'd206;
		10'd632  :  out_col <= 8'd206;
		10'd633  :  out_col <= 8'd206;
		10'd634  :  out_col <= 8'd206;
		10'd635  :  out_col <= 8'd207;
		10'd636  :  out_col <= 8'd207;
		10'd637  :  out_col <= 8'd207;
		10'd638  :  out_col <= 8'd207;
		10'd639  :  out_col <= 8'd207;
		10'd640  :  out_col <= 8'd207;
		10'd641  :  out_col <= 8'd207;
		10'd642  :  out_col <= 8'd208;
		10'd643  :  out_col <= 8'd208;
		10'd644  :  out_col <= 8'd208;
		10'd645  :  out_col <= 8'd208;
		10'd646  :  out_col <= 8'd208;
		10'd647  :  out_col <= 8'd208;
		10'd648  :  out_col <= 8'd208;
		10'd649  :  out_col <= 8'd209;
		10'd650  :  out_col <= 8'd209;
		10'd651  :  out_col <= 8'd209;
		10'd652  :  out_col <= 8'd209;
		10'd653  :  out_col <= 8'd209;
		10'd654  :  out_col <= 8'd209;
		10'd655  :  out_col <= 8'd209;
		10'd656  :  out_col <= 8'd210;
		10'd657  :  out_col <= 8'd210;
		10'd658  :  out_col <= 8'd210;
		10'd659  :  out_col <= 8'd210;
		10'd660  :  out_col <= 8'd210;
		10'd661  :  out_col <= 8'd210;
		10'd662  :  out_col <= 8'd210;
		10'd663  :  out_col <= 8'd211;
		10'd664  :  out_col <= 8'd211;
		10'd665  :  out_col <= 8'd211;
		10'd666  :  out_col <= 8'd211;
		10'd667  :  out_col <= 8'd211;
		10'd668  :  out_col <= 8'd211;
		10'd669  :  out_col <= 8'd211;
		10'd670  :  out_col <= 8'd212;
		10'd671  :  out_col <= 8'd212;
		10'd672  :  out_col <= 8'd212;
		10'd673  :  out_col <= 8'd212;
		10'd674  :  out_col <= 8'd212;
		10'd675  :  out_col <= 8'd212;
		10'd676  :  out_col <= 8'd212;
		10'd677  :  out_col <= 8'd212;
		10'd678  :  out_col <= 8'd213;
		10'd679  :  out_col <= 8'd213;
		10'd680  :  out_col <= 8'd213;
		10'd681  :  out_col <= 8'd213;
		10'd682  :  out_col <= 8'd213;
		10'd683  :  out_col <= 8'd213;
		10'd684  :  out_col <= 8'd213;
		10'd685  :  out_col <= 8'd214;
		10'd686  :  out_col <= 8'd214;
		10'd687  :  out_col <= 8'd214;
		10'd688  :  out_col <= 8'd214;
		10'd689  :  out_col <= 8'd214;
		10'd690  :  out_col <= 8'd214;
		10'd691  :  out_col <= 8'd214;
		10'd692  :  out_col <= 8'd215;
		10'd693  :  out_col <= 8'd215;
		10'd694  :  out_col <= 8'd215;
		10'd695  :  out_col <= 8'd215;
		10'd696  :  out_col <= 8'd215;
		10'd697  :  out_col <= 8'd215;
		10'd698  :  out_col <= 8'd215;
		10'd699  :  out_col <= 8'd216;
		10'd700  :  out_col <= 8'd216;
		10'd701  :  out_col <= 8'd216;
		10'd702  :  out_col <= 8'd216;
		10'd703  :  out_col <= 8'd216;
		10'd704  :  out_col <= 8'd216;
		10'd705  :  out_col <= 8'd216;
		10'd706  :  out_col <= 8'd216;
		10'd707  :  out_col <= 8'd217;
		10'd708  :  out_col <= 8'd217;
		10'd709  :  out_col <= 8'd217;
		10'd710  :  out_col <= 8'd217;
		10'd711  :  out_col <= 8'd217;
		10'd712  :  out_col <= 8'd217;
		10'd713  :  out_col <= 8'd217;
		10'd714  :  out_col <= 8'd218;
		10'd715  :  out_col <= 8'd218;
		10'd716  :  out_col <= 8'd218;
		10'd717  :  out_col <= 8'd218;
		10'd718  :  out_col <= 8'd218;
		10'd719  :  out_col <= 8'd218;
		10'd720  :  out_col <= 8'd218;
		10'd721  :  out_col <= 8'd219;
		10'd722  :  out_col <= 8'd219;
		10'd723  :  out_col <= 8'd219;
		10'd724  :  out_col <= 8'd219;
		10'd725  :  out_col <= 8'd219;
		10'd726  :  out_col <= 8'd219;
		10'd727  :  out_col <= 8'd219;
		10'd728  :  out_col <= 8'd219;
		10'd729  :  out_col <= 8'd220;
		10'd730  :  out_col <= 8'd220;
		10'd731  :  out_col <= 8'd220;
		10'd732  :  out_col <= 8'd220;
		10'd733  :  out_col <= 8'd220;
		10'd734  :  out_col <= 8'd220;
		10'd735  :  out_col <= 8'd220;
		10'd736  :  out_col <= 8'd221;
		10'd737  :  out_col <= 8'd221;
		10'd738  :  out_col <= 8'd221;
		10'd739  :  out_col <= 8'd221;
		10'd740  :  out_col <= 8'd221;
		10'd741  :  out_col <= 8'd221;
		10'd742  :  out_col <= 8'd221;
		10'd743  :  out_col <= 8'd221;
		10'd744  :  out_col <= 8'd222;
		10'd745  :  out_col <= 8'd222;
		10'd746  :  out_col <= 8'd222;
		10'd747  :  out_col <= 8'd222;
		10'd748  :  out_col <= 8'd222;
		10'd749  :  out_col <= 8'd222;
		10'd750  :  out_col <= 8'd222;
		10'd751  :  out_col <= 8'd222;
		10'd752  :  out_col <= 8'd223;
		10'd753  :  out_col <= 8'd223;
		10'd754  :  out_col <= 8'd223;
		10'd755  :  out_col <= 8'd223;
		10'd756  :  out_col <= 8'd223;
		10'd757  :  out_col <= 8'd223;
		10'd758  :  out_col <= 8'd223;
		10'd759  :  out_col <= 8'd224;
		10'd760  :  out_col <= 8'd224;
		10'd761  :  out_col <= 8'd224;
		10'd762  :  out_col <= 8'd224;
		10'd763  :  out_col <= 8'd224;
		10'd764  :  out_col <= 8'd224;
		10'd765  :  out_col <= 8'd224;
		10'd766  :  out_col <= 8'd224;
		10'd767  :  out_col <= 8'd225;
		10'd768  :  out_col <= 8'd225;
		10'd769  :  out_col <= 8'd225;
		10'd770  :  out_col <= 8'd225;
		10'd771  :  out_col <= 8'd225;
		10'd772  :  out_col <= 8'd225;
		10'd773  :  out_col <= 8'd225;
		10'd774  :  out_col <= 8'd225;
		10'd775  :  out_col <= 8'd226;
		10'd776  :  out_col <= 8'd226;
		10'd777  :  out_col <= 8'd226;
		10'd778  :  out_col <= 8'd226;
		10'd779  :  out_col <= 8'd226;
		10'd780  :  out_col <= 8'd226;
		10'd781  :  out_col <= 8'd226;
		10'd782  :  out_col <= 8'd227;
		10'd783  :  out_col <= 8'd227;
		10'd784  :  out_col <= 8'd227;
		10'd785  :  out_col <= 8'd227;
		10'd786  :  out_col <= 8'd227;
		10'd787  :  out_col <= 8'd227;
		10'd788  :  out_col <= 8'd227;
		10'd789  :  out_col <= 8'd227;
		10'd790  :  out_col <= 8'd228;
		10'd791  :  out_col <= 8'd228;
		10'd792  :  out_col <= 8'd228;
		10'd793  :  out_col <= 8'd228;
		10'd794  :  out_col <= 8'd228;
		10'd795  :  out_col <= 8'd228;
		10'd796  :  out_col <= 8'd228;
		10'd797  :  out_col <= 8'd228;
		10'd798  :  out_col <= 8'd229;
		10'd799  :  out_col <= 8'd229;
		10'd800  :  out_col <= 8'd229;
		10'd801  :  out_col <= 8'd229;
		10'd802  :  out_col <= 8'd229;
		10'd803  :  out_col <= 8'd229;
		10'd804  :  out_col <= 8'd229;
		10'd805  :  out_col <= 8'd229;
		10'd806  :  out_col <= 8'd230;
		10'd807  :  out_col <= 8'd230;
		10'd808  :  out_col <= 8'd230;
		10'd809  :  out_col <= 8'd230;
		10'd810  :  out_col <= 8'd230;
		10'd811  :  out_col <= 8'd230;
		10'd812  :  out_col <= 8'd230;
		10'd813  :  out_col <= 8'd230;
		10'd814  :  out_col <= 8'd231;
		10'd815  :  out_col <= 8'd231;
		10'd816  :  out_col <= 8'd231;
		10'd817  :  out_col <= 8'd231;
		10'd818  :  out_col <= 8'd231;
		10'd819  :  out_col <= 8'd231;
		10'd820  :  out_col <= 8'd231;
		10'd821  :  out_col <= 8'd231;
		10'd822  :  out_col <= 8'd232;
		10'd823  :  out_col <= 8'd232;
		10'd824  :  out_col <= 8'd232;
		10'd825  :  out_col <= 8'd232;
		10'd826  :  out_col <= 8'd232;
		10'd827  :  out_col <= 8'd232;
		10'd828  :  out_col <= 8'd232;
		10'd829  :  out_col <= 8'd232;
		10'd830  :  out_col <= 8'd233;
		10'd831  :  out_col <= 8'd233;
		10'd832  :  out_col <= 8'd233;
		10'd833  :  out_col <= 8'd233;
		10'd834  :  out_col <= 8'd233;
		10'd835  :  out_col <= 8'd233;
		10'd836  :  out_col <= 8'd233;
		10'd837  :  out_col <= 8'd233;
		10'd838  :  out_col <= 8'd234;
		10'd839  :  out_col <= 8'd234;
		10'd840  :  out_col <= 8'd234;
		10'd841  :  out_col <= 8'd234;
		10'd842  :  out_col <= 8'd234;
		10'd843  :  out_col <= 8'd234;
		10'd844  :  out_col <= 8'd234;
		10'd845  :  out_col <= 8'd234;
		10'd846  :  out_col <= 8'd235;
		10'd847  :  out_col <= 8'd235;
		10'd848  :  out_col <= 8'd235;
		10'd849  :  out_col <= 8'd235;
		10'd850  :  out_col <= 8'd235;
		10'd851  :  out_col <= 8'd235;
		10'd852  :  out_col <= 8'd235;
		10'd853  :  out_col <= 8'd235;
		10'd854  :  out_col <= 8'd236;
		10'd855  :  out_col <= 8'd236;
		10'd856  :  out_col <= 8'd236;
		10'd857  :  out_col <= 8'd236;
		10'd858  :  out_col <= 8'd236;
		10'd859  :  out_col <= 8'd236;
		10'd860  :  out_col <= 8'd236;
		10'd861  :  out_col <= 8'd236;
		10'd862  :  out_col <= 8'd236;
		10'd863  :  out_col <= 8'd237;
		10'd864  :  out_col <= 8'd237;
		10'd865  :  out_col <= 8'd237;
		10'd866  :  out_col <= 8'd237;
		10'd867  :  out_col <= 8'd237;
		10'd868  :  out_col <= 8'd237;
		10'd869  :  out_col <= 8'd237;
		10'd870  :  out_col <= 8'd237;
		10'd871  :  out_col <= 8'd238;
		10'd872  :  out_col <= 8'd238;
		10'd873  :  out_col <= 8'd238;
		10'd874  :  out_col <= 8'd238;
		10'd875  :  out_col <= 8'd238;
		10'd876  :  out_col <= 8'd238;
		10'd877  :  out_col <= 8'd238;
		10'd878  :  out_col <= 8'd238;
		10'd879  :  out_col <= 8'd239;
		10'd880  :  out_col <= 8'd239;
		10'd881  :  out_col <= 8'd239;
		10'd882  :  out_col <= 8'd239;
		10'd883  :  out_col <= 8'd239;
		10'd884  :  out_col <= 8'd239;
		10'd885  :  out_col <= 8'd239;
		10'd886  :  out_col <= 8'd239;
		10'd887  :  out_col <= 8'd239;
		10'd888  :  out_col <= 8'd240;
		10'd889  :  out_col <= 8'd240;
		10'd890  :  out_col <= 8'd240;
		10'd891  :  out_col <= 8'd240;
		10'd892  :  out_col <= 8'd240;
		10'd893  :  out_col <= 8'd240;
		10'd894  :  out_col <= 8'd240;
		10'd895  :  out_col <= 8'd240;
		10'd896  :  out_col <= 8'd241;
		10'd897  :  out_col <= 8'd241;
		10'd898  :  out_col <= 8'd241;
		10'd899  :  out_col <= 8'd241;
		10'd900  :  out_col <= 8'd241;
		10'd901  :  out_col <= 8'd241;
		10'd902  :  out_col <= 8'd241;
		10'd903  :  out_col <= 8'd241;
		10'd904  :  out_col <= 8'd241;
		10'd905  :  out_col <= 8'd242;
		10'd906  :  out_col <= 8'd242;
		10'd907  :  out_col <= 8'd242;
		10'd908  :  out_col <= 8'd242;
		10'd909  :  out_col <= 8'd242;
		10'd910  :  out_col <= 8'd242;
		10'd911  :  out_col <= 8'd242;
		10'd912  :  out_col <= 8'd242;
		10'd913  :  out_col <= 8'd243;
		10'd914  :  out_col <= 8'd243;
		10'd915  :  out_col <= 8'd243;
		10'd916  :  out_col <= 8'd243;
		10'd917  :  out_col <= 8'd243;
		10'd918  :  out_col <= 8'd243;
		10'd919  :  out_col <= 8'd243;
		10'd920  :  out_col <= 8'd243;
		10'd921  :  out_col <= 8'd243;
		10'd922  :  out_col <= 8'd244;
		10'd923  :  out_col <= 8'd244;
		10'd924  :  out_col <= 8'd244;
		10'd925  :  out_col <= 8'd244;
		10'd926  :  out_col <= 8'd244;
		10'd927  :  out_col <= 8'd244;
		10'd928  :  out_col <= 8'd244;
		10'd929  :  out_col <= 8'd244;
		10'd930  :  out_col <= 8'd245;
		10'd931  :  out_col <= 8'd245;
		10'd932  :  out_col <= 8'd245;
		10'd933  :  out_col <= 8'd245;
		10'd934  :  out_col <= 8'd245;
		10'd935  :  out_col <= 8'd245;
		10'd936  :  out_col <= 8'd245;
		10'd937  :  out_col <= 8'd245;
		10'd938  :  out_col <= 8'd245;
		10'd939  :  out_col <= 8'd246;
		10'd940  :  out_col <= 8'd246;
		10'd941  :  out_col <= 8'd246;
		10'd942  :  out_col <= 8'd246;
		10'd943  :  out_col <= 8'd246;
		10'd944  :  out_col <= 8'd246;
		10'd945  :  out_col <= 8'd246;
		10'd946  :  out_col <= 8'd246;
		10'd947  :  out_col <= 8'd246;
		10'd948  :  out_col <= 8'd247;
		10'd949  :  out_col <= 8'd247;
		10'd950  :  out_col <= 8'd247;
		10'd951  :  out_col <= 8'd247;
		10'd952  :  out_col <= 8'd247;
		10'd953  :  out_col <= 8'd247;
		10'd954  :  out_col <= 8'd247;
		10'd955  :  out_col <= 8'd247;
		10'd956  :  out_col <= 8'd248;
		10'd957  :  out_col <= 8'd248;
		10'd958  :  out_col <= 8'd248;
		10'd959  :  out_col <= 8'd248;
		10'd960  :  out_col <= 8'd248;
		10'd961  :  out_col <= 8'd248;
		10'd962  :  out_col <= 8'd248;
		10'd963  :  out_col <= 8'd248;
		10'd964  :  out_col <= 8'd248;
		10'd965  :  out_col <= 8'd249;
		10'd966  :  out_col <= 8'd249;
		10'd967  :  out_col <= 8'd249;
		10'd968  :  out_col <= 8'd249;
		10'd969  :  out_col <= 8'd249;
		10'd970  :  out_col <= 8'd249;
		10'd971  :  out_col <= 8'd249;
		10'd972  :  out_col <= 8'd249;
		10'd973  :  out_col <= 8'd249;
		10'd974  :  out_col <= 8'd250;
		10'd975  :  out_col <= 8'd250;
		10'd976  :  out_col <= 8'd250;
		10'd977  :  out_col <= 8'd250;
		10'd978  :  out_col <= 8'd250;
		10'd979  :  out_col <= 8'd250;
		10'd980  :  out_col <= 8'd250;
		10'd981  :  out_col <= 8'd250;
		10'd982  :  out_col <= 8'd250;
		10'd983  :  out_col <= 8'd251;
		10'd984  :  out_col <= 8'd251;
		10'd985  :  out_col <= 8'd251;
		10'd986  :  out_col <= 8'd251;
		10'd987  :  out_col <= 8'd251;
		10'd988  :  out_col <= 8'd251;
		10'd989  :  out_col <= 8'd251;
		10'd990  :  out_col <= 8'd251;
		10'd991  :  out_col <= 8'd251;
		10'd992  :  out_col <= 8'd252;
		10'd993  :  out_col <= 8'd252;
		10'd994  :  out_col <= 8'd252;
		10'd995  :  out_col <= 8'd252;
		10'd996  :  out_col <= 8'd252;
		10'd997  :  out_col <= 8'd252;
		10'd998  :  out_col <= 8'd252;
		10'd999  :  out_col <= 8'd252;
		10'd1000  :  out_col <= 8'd252;
		10'd1001  :  out_col <= 8'd253;
		10'd1002  :  out_col <= 8'd253;
		10'd1003  :  out_col <= 8'd253;
		10'd1004  :  out_col <= 8'd253;
		10'd1005  :  out_col <= 8'd253;
		10'd1006  :  out_col <= 8'd253;
		10'd1007  :  out_col <= 8'd253;
		10'd1008  :  out_col <= 8'd253;
		10'd1009  :  out_col <= 8'd253;
		10'd1010  :  out_col <= 8'd254;
		10'd1011  :  out_col <= 8'd254;
		10'd1012  :  out_col <= 8'd254;
		10'd1013  :  out_col <= 8'd254;
		10'd1014  :  out_col <= 8'd254;
		10'd1015  :  out_col <= 8'd254;
		10'd1016  :  out_col <= 8'd254;
		10'd1017  :  out_col <= 8'd254;
		10'd1018  :  out_col <= 8'd254;
		10'd1019  :  out_col <= 8'd255;
		10'd1020  :  out_col <= 8'd255;
		10'd1021  :  out_col <= 8'd255;
		10'd1022  :  out_col <= 8'd255;
		10'd1023  :  out_col <= 8'd255;
		default   :  out_col <= 8'd0;
	endcase
end
endmodule
